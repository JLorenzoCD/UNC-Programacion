`timescale 1ns / 1ps

module execute_tb;

endmodule
